`define NOERROR         2'b00
`define RXSTARTERROR    2'b01
`define RXPARITYERROR   2'b10
`define RXSTOPERROR     2'b11
