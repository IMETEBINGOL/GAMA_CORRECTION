// Generated Verilog Header File
// This file is automatically generated from an Excel file.

RandomAccessMemory[0] <= 16'd266;
RandomAccessMemory[1] <= 16'd0;
RandomAccessMemory[2] <= 16'd0;
RandomAccessMemory[3] <= 16'd0;
RandomAccessMemory[4] <= 16'd0;
RandomAccessMemory[5] <= 16'd0;
RandomAccessMemory[6] <= 16'd0;
RandomAccessMemory[7] <= 16'd0;
RandomAccessMemory[8] <= 16'd0;
RandomAccessMemory[9] <= 16'd0;
RandomAccessMemory[10] <= 16'd0;
RandomAccessMemory[11] <= 16'd0;
RandomAccessMemory[12] <= 16'd0;
RandomAccessMemory[13] <= 16'd0;
RandomAccessMemory[14] <= 16'd0;
RandomAccessMemory[15] <= 16'd0;
RandomAccessMemory[16] <= 16'd0;
RandomAccessMemory[17] <= 16'd0;
RandomAccessMemory[18] <= 16'd0;
RandomAccessMemory[19] <= 16'd0;
RandomAccessMemory[20] <= 16'd0;
RandomAccessMemory[21] <= 16'd0;
RandomAccessMemory[22] <= 16'd0;
RandomAccessMemory[23] <= 16'd0;
RandomAccessMemory[24] <= 16'd0;
RandomAccessMemory[25] <= 16'd0;
RandomAccessMemory[26] <= 16'd0;
RandomAccessMemory[27] <= 16'd0;
RandomAccessMemory[28] <= 16'd0;
RandomAccessMemory[29] <= 16'd0;
RandomAccessMemory[30] <= 16'd0;
RandomAccessMemory[31] <= 16'd0;
RandomAccessMemory[32] <= 16'd0;
RandomAccessMemory[33] <= 16'd0;
RandomAccessMemory[34] <= 16'd0;
RandomAccessMemory[35] <= 16'd0;
RandomAccessMemory[36] <= 16'd0;
RandomAccessMemory[37] <= 16'd0;
RandomAccessMemory[38] <= 16'd0;
RandomAccessMemory[39] <= 16'd0;
RandomAccessMemory[40] <= 16'd0;
RandomAccessMemory[41] <= 16'd0;
RandomAccessMemory[42] <= 16'd0;
RandomAccessMemory[43] <= 16'd0;
RandomAccessMemory[44] <= 16'd0;
RandomAccessMemory[45] <= 16'd0;
RandomAccessMemory[46] <= 16'd0;
RandomAccessMemory[47] <= 16'd0;
RandomAccessMemory[48] <= 16'd0;
RandomAccessMemory[49] <= 16'd0;
RandomAccessMemory[50] <= 16'd0;
RandomAccessMemory[51] <= 16'd0;
RandomAccessMemory[52] <= 16'd0;
RandomAccessMemory[53] <= 16'd0;
RandomAccessMemory[54] <= 16'd0;
RandomAccessMemory[55] <= 16'd0;
RandomAccessMemory[56] <= 16'd0;
RandomAccessMemory[57] <= 16'd0;
RandomAccessMemory[58] <= 16'd0;
RandomAccessMemory[59] <= 16'd0;
RandomAccessMemory[60] <= 16'd0;
RandomAccessMemory[61] <= 16'd0;
RandomAccessMemory[62] <= 16'd0;
RandomAccessMemory[63] <= 16'd0;
RandomAccessMemory[64] <= 16'd0;
RandomAccessMemory[65] <= 16'd0;
RandomAccessMemory[66] <= 16'd0;
RandomAccessMemory[67] <= 16'd0;
RandomAccessMemory[68] <= 16'd0;
RandomAccessMemory[69] <= 16'd0;
RandomAccessMemory[70] <= 16'd0;
RandomAccessMemory[71] <= 16'd0;
RandomAccessMemory[72] <= 16'd0;
RandomAccessMemory[73] <= 16'd0;
RandomAccessMemory[74] <= 16'd0;
RandomAccessMemory[75] <= 16'd0;
RandomAccessMemory[76] <= 16'd0;
RandomAccessMemory[77] <= 16'd0;
RandomAccessMemory[78] <= 16'd0;
RandomAccessMemory[79] <= 16'd0;
RandomAccessMemory[80] <= 16'd0;
RandomAccessMemory[81] <= 16'd0;
RandomAccessMemory[82] <= 16'd0;
RandomAccessMemory[83] <= 16'd0;
RandomAccessMemory[84] <= 16'd0;
RandomAccessMemory[85] <= 16'd0;
RandomAccessMemory[86] <= 16'd0;
RandomAccessMemory[87] <= 16'd0;
RandomAccessMemory[88] <= 16'd0;
RandomAccessMemory[89] <= 16'd0;
RandomAccessMemory[90] <= 16'd0;
RandomAccessMemory[91] <= 16'd0;
RandomAccessMemory[92] <= 16'd0;
RandomAccessMemory[93] <= 16'd0;
RandomAccessMemory[94] <= 16'd0;
RandomAccessMemory[95] <= 16'd0;
RandomAccessMemory[96] <= 16'd0;
RandomAccessMemory[97] <= 16'd0;
RandomAccessMemory[98] <= 16'd0;
RandomAccessMemory[99] <= 16'd0;
RandomAccessMemory[100] <= 16'd0;
RandomAccessMemory[101] <= 16'd0;
RandomAccessMemory[102] <= 16'd0;
RandomAccessMemory[103] <= 16'd0;
RandomAccessMemory[104] <= 16'd0;
RandomAccessMemory[105] <= 16'd0;
RandomAccessMemory[106] <= 16'd0;
RandomAccessMemory[107] <= 16'd0;
RandomAccessMemory[108] <= 16'd0;
RandomAccessMemory[109] <= 16'd0;
RandomAccessMemory[110] <= 16'd0;
RandomAccessMemory[111] <= 16'd0;
RandomAccessMemory[112] <= 16'd0;
RandomAccessMemory[113] <= 16'd0;
RandomAccessMemory[114] <= 16'd0;
RandomAccessMemory[115] <= 16'd0;
RandomAccessMemory[116] <= 16'd0;
RandomAccessMemory[117] <= 16'd0;
RandomAccessMemory[118] <= 16'd0;
RandomAccessMemory[119] <= 16'd0;
RandomAccessMemory[120] <= 16'd0;
RandomAccessMemory[121] <= 16'd0;
RandomAccessMemory[122] <= 16'd0;
RandomAccessMemory[123] <= 16'd0;
RandomAccessMemory[124] <= 16'd0;
RandomAccessMemory[125] <= 16'd0;
RandomAccessMemory[126] <= 16'd0;
RandomAccessMemory[127] <= 16'd0;
