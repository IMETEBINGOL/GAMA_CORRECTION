default:
begin
    resetState;
end