`define getUartErrorOpcode      8'h01
`define readSettingsOpcode      8'h02
`define resetFifoOpcode         8'h03
`define resetSettingsOpcode     8'h04
`define writeSettingsOpcode     8'h05
